package tb_tasks;

task Seg_initial(input clk);
	
endtask : Seg_initial

endpackage : tb_tasks