package tb_tasks;
	
task Seg_initial();
	
endtask : Seg_initial
endpackage : tb_tasks