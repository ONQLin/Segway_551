`define TP2